`include "ral_reg_block.sv"

`include "ral_adapter.sv"

`include "ral_sequence.sv"

`include "ral_sequencer.sv"

`include "ral_driver.sv"

`include "ral_monitor.sv"

`include "ral_scoreboard.sv"

`include "ral_agent.sv"

`include "ral_env.sv"

`include "ral_test.sv"

 
