
package ral_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ral_reg_ctrl.sv"
  `include "ral_reg_Reg1.sv"
  `include "ral_reg_Reg2.sv"
  `include "ral_reg_Reg3.sv"
  `include "ral_reg_Reg4.sv"
  `include "ral_block.sv"

endpackage
